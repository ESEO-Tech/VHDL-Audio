
package OscillatorTestbench_pkg is
	constant CLK_FREQUENCY_HZ   : positive := 51_200_000;
	constant OSC_SAMPLE_RATE_HZ : positive := 20_000;
    constant OSC_STEP           : positive := 7;
end OscillatorTestbench_pkg;
