
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity I2STransmitter is
	generic (
        -- Generic parameter declarations.
	);
	port (
        -- Port declarations.
	);
end I2STransmitter;

architecture RTL of I2STransmitter is
    -- Type, constant and signal declarations.
begin
    -- Concurrent statements.
end RTL;
